../../ODMB/LED_ODMB7/TEST/LED_test_v2/LED_test_v2.srcs/sources_1/imports/new/LED_blinker.vhd